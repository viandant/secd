

-- Automatically generated SECD microcode

library ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity microcode_rom is
  port (clk  : in std_logic;
        en   : in std_logic;
        addr : in std_logic_vector(8 downto 0);
        data : out std_logic_vector(27 downto 0));
end microcode_rom;

architecture rtl of microcode_rom is

constant MICROCODE_ROM_SIZE : integer := 512;
type rom_type is array (0 to MICROCODE_ROM_SIZE - 1) of std_logic_vector (27 downto 0);
constant MICROCODE_ROM : rom_type := (
"0000101110001000000000000000", -- 0                                                         jump      boot
"0001100000001000000000000000", -- 1   ld-ins                                                jump      ld
"0010101110001000000000000000", -- 2   ldc-ins                                               jump      ldc
"0011000100001000000000000000", -- 3   ldf-ins                                               jump      ldf
"0011011110001000000000000000", -- 4   ap-ins                                                jump      ap
"0100010110001000000000000000", -- 5   rtn-ins                                               jump      rtn
"0100111100001000000000000000", -- 6   dum-ins                                               jump      dum
"0101000110001000000000000000", -- 7   rap-ins                                               jump      rap
"0110000100001000000000000000", -- 8   sel-ins                                               jump      sel
"0110111100001000000000000000", -- 9   join-ins                                              jump      join
"0111001000001000000000000000", -- 10  car-ins                                               jump      car
"0111011100001000000000000000", -- 11  cdr-ins                                               jump      cdr
"0111101110001000000000000000", -- 12  atom-ins                                              jump      atom
"1000000100001000000000000000", -- 13  cons-ins                                              jump      cons
"1000100100001000000000000000", -- 14  eq-ins                                                jump      eq
"1000110000001000000000000000", -- 15  add-ins                                               jump      add
"1000111000001000000000000000", -- 16  sub-ins                                               jump      sub
"1001000000001000000000000000", -- 17  mul-ins                                               jump      mul
"1001001000001000000000000000", -- 18  div-ins                                               jump      div
"1001010000001000000000000000", -- 19  rem-ins                                               jump      rem
"1001011000001000000000000000", -- 20  leq-ins                                               jump      leq
"1001100100001000000000000000", -- 21  stop-ins                                              jump      stop
"1001101110001000000000000000", -- 22  external-ins                                          jump      external
"0000111011011100010000000000", -- 23  boot            1                         halted      button?   start-program
"0000101110001000000000000000", -- 24                                                        jump      boot
"0000110111011000000000000000", -- 25  error           2                                     button?   _3
"0000110010001000000000000000", -- 26                                                        jump      error
"0000110111011000000000000000", -- 27  _3                                                    button?   _3
"0000101110001000000000000000", -- 28                                                        jump      boot
"0000000000000100000101010011", -- 29  start-program       num        mar        running     
"0000000000000000000010100010", -- 30                      mem        car                    
"0000000000000000000101000110", -- 31                      car        mar                    
"0000000000000000000011000010", -- 32                      mem        s                      
"0000000000000000000011110100", -- 33                      nilx       e                      
"0000000000000000000101010011", -- 34                      num        mar                    
"0000000000000000000010100010", -- 35                      mem        car                    
"0000000000000000000101000110", -- 36                      car        mar                    
"0000000000000000000010100010", -- 37                      mem        car                    
"0000000000000000000100000110", -- 38                      car        c                      
"0000000000000000000100110100", -- 39                      nilx       d                      
"0000000000000000000101110100", -- 40                      nilx       x1                     
"0000000000000000000110010100", -- 41                      nilx       x2                     
"0000000000000000000101010011", -- 42                      num        mar                    
"0000000000000000000110100010", -- 43                      mem        free                   
"0000000000000000000101001001", -- 44  top-of-cycle        c          mar                    
"0000000000000000000010100010", -- 45                      mem        car                    
"0000000000000000000101000110", -- 46                      car        mar                    
"0000000000010000000001000010", -- 47                      mem        arg                    dispatch  
"0000000000000000000101101000", -- 48  ld                  e          x1                     
"0000000000000000000101001001", -- 49                      c          mar                    
"0000000000000000000110000010", -- 50                      mem        x2                     
"0000000000000000000101001101", -- 51                      x2         mar                    
"0000000000000000000010100010", -- 52                      mem        car                    
"0000000000000000000101000110", -- 53                      car        mar                    
"0000000000000000000010100010", -- 54                      mem        car                    
"0000000000000000000101000110", -- 55                      car        mar                    
"0000000000000000000001000010", -- 56                      mem        arg                    
"0001111101010000000000000011", -- 57  _7                  arg                               nil?      _8
"0000000000000000000101001100", -- 58                      x1         mar                    
"0000000000000000000101100010", -- 59                      mem        x1                     
"0000000000000000010001100000", -- 60                                 buf1       dec         
"0001110010001000000001000100", -- 61                      buf1       arg                    jump      _7
"0000000000000000000101001100", -- 62  _8                  x1         mar                    
"0000000000000000000010100010", -- 63                      mem        car                    
"0000000000000000000101100110", -- 64                      car        x1                     
"0000000000000000000101001001", -- 65                      c          mar                    
"0000000000000000000110000010", -- 66                      mem        x2                     
"0000000000000000000101001101", -- 67                      x2         mar                    
"0000000000000000000010100010", -- 68                      mem        car                    
"0000000000000000000101000110", -- 69                      car        mar                    
"0000000000000000000110000010", -- 70                      mem        x2                     
"0000000000000000000101001101", -- 71                      x2         mar                    
"0000000000000000000001000010", -- 72                      mem        arg                    
"0010011101010000000000000011", -- 73  _9                  arg                               nil?      _10
"0000000000000000000101001100", -- 74                      x1         mar                    
"0000000000000000000101100010", -- 75                      mem        x1                     
"0000000000000000010001100000", -- 76                                 buf1       dec         
"0010010010001000000001000100", -- 77                      buf1       arg                    jump      _9
"0000000000000000000101001100", -- 78  _10                 x1         mar                    
"0000000000000000000010100010", -- 79                      mem        car                    
"0000000000000000000101100110", -- 80                      car        x1                     
"1010010111100000000110000111", -- 81                      s          x2                     call      consx1x2
"0000000000000000000011001011", -- 82                      mar        s                      
"0000000000000000000101001001", -- 83                      c          mar                    
"0000000000000000000100000010", -- 84                      mem        c                      
"0000000000000000000101001001", -- 85                      c          mar                    
"0001011000001000000100000010", -- 86                      mem        c                      jump      top-of-cycle
"0000000000000000000110000111", -- 87  ldc                 s          x2                     
"0000000000000000000101001001", -- 88                      c          mar                    
"0000000000000000000101100010", -- 89                      mem        x1                     
"0000000000000000000101001100", -- 90                      x1         mar                    
"0000000000000000000010100010", -- 91                      mem        car                    
"1010010111100000000101100110", -- 92                      car        x1                     call      consx1x2
"0000000000000000000011001011", -- 93                      mar        s                      
"0000000000000000000101001001", -- 94                      c          mar                    
"0000000000000000000100000010", -- 95                      mem        c                      
"0000000000000000000101001001", -- 96                      c          mar                    
"0001011000001000000100000010", -- 97                      mem        c                      jump      top-of-cycle
"0000000000000000000110001000", -- 98  ldf                 e          x2                     
"0000000000000000000101001001", -- 99                      c          mar                    
"0000000000000000000101100010", -- 100                     mem        x1                     
"0000000000000000000101001100", -- 101                     x1         mar                    
"0000000000000000000010100010", -- 102                     mem        car                    
"1010010111100000000101100110", -- 103                     car        x1                     call      consx1x2
"0000000000000000000101101011", -- 104                     mar        x1                     
"1010010111100000000110000111", -- 105                     s          x2                     call      consx1x2
"0000000000000000000011001011", -- 106                     mar        s                      
"0000000000000000000101001001", -- 107                     c          mar                    
"0000000000000000000100000010", -- 108                     mem        c                      
"0000000000000000000101001001", -- 109                     c          mar                    
"0001011000001000000100000010", -- 110                     mem        c                      jump      top-of-cycle
"0000000000000000000110001010", -- 111 ap                  d          x2                     
"0000000000000000000101001001", -- 112                     c          mar                    
"1010010111100000000101100010", -- 113                     mem        x1                     call      consx1x2
"0000000000000000000110001011", -- 114                     mar        x2                     
"1010010111100000000101101000", -- 115                     e          x1                     call      consx1x2
"0000000000000000000110001011", -- 116                     mar        x2                     
"0000000000000000000101000111", -- 117                     s          mar                    
"0000000000000000000101100010", -- 118                     mem        x1                     
"0000000000000000000101001100", -- 119                     x1         mar                    
"1010010111100000000101100010", -- 120                     mem        x1                     call      consx1x2
"0000000000000000000100101011", -- 121                     mar        d                      
"0000000000000000000101000111", -- 122                     s          mar                    
"0000000000000000000010100010", -- 123                     mem        car                    
"0000000000000000000101000110", -- 124                     car        mar                    
"0000000000000000000110000010", -- 125                     mem        x2                     
"0000000000000000000101000111", -- 126                     s          mar                    
"0000000000000000000101100010", -- 127                     mem        x1                     
"0000000000000000000101001100", -- 128                     x1         mar                    
"0000000000000000000010100010", -- 129                     mem        car                    
"1010010111100000000101100110", -- 130                     car        x1                     call      consx1x2
"0000000000000000000011101011", -- 131                     mar        e                      
"0000000000000000000000000000", -- 132                                                       
"0000000000000000000101000111", -- 133                     s          mar                    
"0000000000000000000010100010", -- 134                     mem        car                    
"0000000000000000000101000110", -- 135                     car        mar                    
"0000000000000000000010100010", -- 136                     mem        car                    
"0000000000000000000100000110", -- 137                     car        c                      
"0001011000001000000011010100", -- 138                     nilx       s                      jump      top-of-cycle
"0000000000000000000101001010", -- 139 rtn                 d          mar                    
"0000000000000000000010100010", -- 140                     mem        car                    
"0000000000000000000110000110", -- 141                     car        x2                     
"0000000000000000000101000111", -- 142                     s          mar                    
"0000000000000000000010100010", -- 143                     mem        car                    
"1010010111100000000101100110", -- 144                     car        x1                     call      consx1x2
"0000000000000000000011001011", -- 145                     mar        s                      
"0000000000000000000101001010", -- 146                     d          mar                    
"0000000000000000000100100010", -- 147                     mem        d                      
"0000000000000000000101001010", -- 148                     d          mar                    
"0000000000000000000010100010", -- 149                     mem        car                    
"0000000000000000000011100110", -- 150                     car        e                      
"0000000000000000000101001010", -- 151                     d          mar                    
"0000000000000000000100100010", -- 152                     mem        d                      
"0000000000000000000101001010", -- 153                     d          mar                    
"0000000000000000000010100010", -- 154                     mem        car                    
"0000000000000000000100000110", -- 155                     car        c                      
"0000000000000000000101001010", -- 156                     d          mar                    
"0001011000001000000100100010", -- 157                     mem        d                      jump      top-of-cycle
"0000000000000000000110001000", -- 158 dum                 e          x2                     
"1010010111100000000101110100", -- 159                     nilx       x1                     call      consx1x2
"0000000000000000000011101011", -- 160                     mar        e                      
"0000000000000000000101001001", -- 161                     c          mar                    
"0001011000001000000100000010", -- 162                     mem        c                      jump      top-of-cycle
"0000000000000000000110001010", -- 163 rap                 d          x2                     
"0000000000000000000101001001", -- 164                     c          mar                    
"1010010111100000000101100010", -- 165                     mem        x1                     call      consx1x2
"0000000000000000000110001011", -- 166                     mar        x2                     
"0000000000000000000101001000", -- 167                     e          mar                    
"1010010111100000000101100010", -- 168                     mem        x1                     call      consx1x2
"0000000000000000000110001011", -- 169                     mar        x2                     
"0000000000000000000101000111", -- 170                     s          mar                    
"0000000000000000000101100010", -- 171                     mem        x1                     
"0000000000000000000101001100", -- 172                     x1         mar                    
"1010010111100000000101100010", -- 173                     mem        x1                     call      consx1x2
"0000000000000000000100101011", -- 174                     mar        d                      
"0000000000000000000101000111", -- 175                     s          mar                    
"0000000000000000000010100010", -- 176                     mem        car                    
"0000000000000000000101000110", -- 177                     car        mar                    
"0000000000000000000011100010", -- 178                     mem        e                      
"0000000000000000000101000111", -- 179                     s          mar                    
"0000000000000000001000100010", -- 180                     mem        y2                     
"0000000000000000000101010010", -- 181                     y2         mar                    
"0000000000000000000010100010", -- 182                     mem        car                    
"0000000000000000001000100110", -- 183                     car        y2                     
"0000000000000000000101001000", -- 184                     e          mar                    
"0000000000000000000001000010", -- 185                     mem        arg                    
"0000000000000010100001100000", -- 186                                buf1       replcar     
"0000000000000000000000100100", -- 187                     buf1       bidir                  
"0000000000000000000101000111", -- 188                     s          mar                    
"0000000000000000000010100010", -- 189                     mem        car                    
"0000000000000000000101000110", -- 190                     car        mar                    
"0000000000000000000010100010", -- 191                     mem        car                    
"0000000000000000000100000110", -- 192                     car        c                      
"0001011000001000000011010100", -- 193                     nilx       s                      jump      top-of-cycle
"0000000000000000000110001010", -- 194 sel                 d          x2                     
"0000000000000000000101001001", -- 195                     c          mar                    
"0000000000000000000101100010", -- 196                     mem        x1                     
"0000000000000000000101001100", -- 197                     x1         mar                    
"0000000000000000000101100010", -- 198                     mem        x1                     
"0000000000000000000101001100", -- 199                     x1         mar                    
"1010010111100000000101100010", -- 200                     mem        x1                     call      consx1x2
"0000000000000000000100101011", -- 201                     mar        d                      
"0000000000000000000101000111", -- 202                     s          mar                    
"0000000000000000000010100010", -- 203                     mem        car                    
"0000000000000000000101000110", -- 204                     car        mar                    
"0000000000000000000001000010", -- 205                     mem        arg                    
"0000000000000000000101010101", -- 206                     true       mar                    
"0110101110110000000000000010", -- 207                     mem                               eq?       _18
"0000000000000000000101001001", -- 208                     c          mar                    
"0000000000000000000100000010", -- 209                     mem        c                      
"0000000000000000000101001001", -- 210                     c          mar                    
"0000000000000000000100000010", -- 211                     mem        c                      
"0000000000000000000101001001", -- 212                     c          mar                    
"0000000000000000000010100010", -- 213                     mem        car                    
"0110111000001000000100000110", -- 214                     car        c                      jump      _19
"0000000000000000000101001001", -- 215 _18                 c          mar                    
"0000000000000000000100000010", -- 216                     mem        c                      
"0000000000000000000101001001", -- 217                     c          mar                    
"0000000000000000000010100010", -- 218                     mem        car                    
"0000000000000000000100000110", -- 219                     car        c                      
"0000000000000000000101000111", -- 220 _19                 s          mar                    
"0001011000001000000011000010", -- 221                     mem        s                      jump      top-of-cycle
"0000000000000000000100001010", -- 222 join                d          c                      
"0000000000000000000101001001", -- 223                     c          mar                    
"0000000000000000000010100010", -- 224                     mem        car                    
"0000000000000000000100000110", -- 225                     car        c                      
"0000000000000000000101001010", -- 226                     d          mar                    
"0001011000001000000100100010", -- 227                     mem        d                      jump      top-of-cycle
"0000000000000000000101000111", -- 228 car                 s          mar                    
"0000000000000000000110000010", -- 229                     mem        x2                     
"0000000000000000000101000111", -- 230                     s          mar                    
"0000000000000000000010100010", -- 231                     mem        car                    
"0000000000000000000101000110", -- 232                     car        mar                    
"0000000000000000000010100010", -- 233                     mem        car                    
"1010010111100000000101100110", -- 234                     car        x1                     call      consx1x2
"0000000000000000000011001011", -- 235                     mar        s                      
"0000000000000000000101001001", -- 236                     c          mar                    
"0001011000001000000100000010", -- 237                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 238 cdr                 s          mar                    
"0000000000000000000110000010", -- 239                     mem        x2                     
"0000000000000000000101000111", -- 240                     s          mar                    
"0000000000000000000010100010", -- 241                     mem        car                    
"0000000000000000000101000110", -- 242                     car        mar                    
"1010010111100000000101100010", -- 243                     mem        x1                     call      consx1x2
"0000000000000000000011001011", -- 244                     mar        s                      
"0000000000000000000101001001", -- 245                     c          mar                    
"0001011000001000000100000010", -- 246                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 247 atom                s          mar                    
"0000000000000000000010100010", -- 248                     mem        car                    
"0000000000000000000101000110", -- 249                     car        mar                    
"0111111001001000000000000010", -- 250                     mem                               atom?     _24
"0111111010001000000101110110", -- 251                     false      x1                     jump      _25
"0000000000000000000101110101", -- 252 _24                 true       x1                     
"0000000000000000000101000111", -- 253 _25                 s          mar                    
"1010010111100000000110000010", -- 254                     mem        x2                     call      consx1x2
"0000000000000000000011001011", -- 255                     mar        s                      
"0000000000000000000101001001", -- 256                     c          mar                    
"0001011000001000000100000010", -- 257                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 258 cons                s          mar                    
"0000000000000000000110000010", -- 259                     mem        x2                     
"0000000000000000000101001101", -- 260                     x2         mar                    
"0000000000000000000010100010", -- 261                     mem        car                    
"0000000000000000000110000110", -- 262                     car        x2                     
"0000000000000000000101000111", -- 263                     s          mar                    
"0000000000000000000010100010", -- 264                     mem        car                    
"1010010111100000000101100110", -- 265                     car        x1                     call      consx1x2
"0000000000000000000101101011", -- 266                     mar        x1                     
"0000000000000000000101000111", -- 267                     s          mar                    
"0000000000000000000110000010", -- 268                     mem        x2                     
"0000000000000000000101001101", -- 269                     x2         mar                    
"1010010111100000000110000010", -- 270                     mem        x2                     call      consx1x2
"0000000000000000000011001011", -- 271                     mar        s                      
"0000000000000000000101001001", -- 272                     c          mar                    
"0001011000001000000100000010", -- 273                     mem        c                      jump      top-of-cycle
"1001110111100000000000000000", -- 274 eq                                                    call      setup-alu-args
"1000101010110000000000000010", -- 275                     mem                               eq?       _28
"1000101100001000000101110110", -- 276                     false      x1                     jump      _29
"0000000000000000000101110101", -- 277 _28                 true       x1                     
"1010001001100000000000000000", -- 278 _29                                                   call      push-alu-result
"0001011000001000000000000000", -- 279                                                       jump      top-of-cycle
"1001110111100000000000000000", -- 280 add                                                   call      setup-alu-args
"1010100011100000100001100010", -- 281                     mem        buf1       add         call      alu-gc
"1010001001100000000101101011", -- 282                     mar        x1                     call      push-alu-result
"0001011000001000000000000000", -- 283                                                       jump      top-of-cycle
"1001110111100000000000000000", -- 284 sub                                                   call      setup-alu-args
"1010100011100000110001100010", -- 285                     mem        buf1       sub         call      alu-gc
"1010001001100000000101101011", -- 286                     mar        x1                     call      push-alu-result
"0001011000001000000000000000", -- 287                                                       jump      top-of-cycle
"1001110111100000000000000000", -- 288 mul                                                   call      setup-alu-args
"1010100011100001000001100010", -- 289                     mem        buf1       mul         call      alu-gc
"1010001001100000000101101011", -- 290                     mar        x1                     call      push-alu-result
"0001011000001000000000000000", -- 291                                                       jump      top-of-cycle
"1001110111100000000000000000", -- 292 div                                                   call      setup-alu-args
"1010100011100001010001100010", -- 293                     mem        buf1       div         call      alu-gc
"1010001001100000000101101011", -- 294                     mar        x1                     call      push-alu-result
"0001011000001000000000000000", -- 295                                                       jump      top-of-cycle
"1001110111100000000000000000", -- 296 rem                                                   call      setup-alu-args
"1010100011100001100001100010", -- 297                     mem        buf1       rem         call      alu-gc
"1010001001100000000101101011", -- 298                     mar        x1                     call      push-alu-result
"0001011000001000000000000000", -- 299                                                       jump      top-of-cycle
"1001110111100000000000000000", -- 300 leq                                                   call      setup-alu-args
"1001011110111000000000000010", -- 301                     mem                               leq?      _36
"1001100000001000000101110110", -- 302                     false      x1                     jump      _37
"0000000000000000000101110101", -- 303 _36                 true       x1                     
"1010001001100000000000000000", -- 304 _37                                                   call      push-alu-result
"0001011000001000000000000000", -- 305                                                       jump      top-of-cycle
"0000000000000000000101000111", -- 306 stop                s          mar                    
"0000000000000000000010100010", -- 307                     mem        car                    
"0000000000000000000011000110", -- 308                     car        s                      
"0000000000000000000101010011", -- 309                     num        mar                    
"0000000001110000000000100111", -- 310                     s          bidir                  stop      
"1001110011011100110000000000", -- 311 external                                  external    button?   external-finish
"1001101110001000000000000000", -- 312                                                       jump      external
"0000000000000100000101001001", -- 313 external-finish     c          mar        running     
"0001011000001000000100000010", -- 314                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 315 setup-alu-args      s          mar                    
"0000000000000000000101100010", -- 316                     mem        x1                     
"0000000000000000000101001100", -- 317                     x1         mar                    
"0000000000000000000010100010", -- 318                     mem        car                    
"0000000000000000000101000110", -- 319                     car        mar                    
"0000000000000000000001000010", -- 320                     mem        arg                    
"0000000000000000000101000111", -- 321                     s          mar                    
"0000000000000000000010100010", -- 322                     mem        car                    
"0000000001101000000101000110", -- 323                     car        mar                    return    
"0000000000000000000101000111", -- 324 push-alu-result     s          mar                    
"0000000000000000000110000010", -- 325                     mem        x2                     
"0000000000000000000101001101", -- 326                     x2         mar                    
"1010010111100000000110000010", -- 327                     mem        x2                     call      consx1x2
"0000000000000000000011001011", -- 328                     mar        s                      
"0000000000000000000101001001", -- 329                     c          mar                    
"0000000001101000000100000010", -- 330                     mem        c                      return    
"1010011111000000000000001110", -- 331 consx1x2            free                              num?      cons-gc
"0000000000000000000101001110", -- 332 _42                 free       mar                    
"0000000000000000000110100010", -- 333                     mem        free                   
"0000000001101000000000110111", -- 334                     cons       bidir                  return    
"1010101111100000000000000000", -- 335 cons-gc                                               call      gc
"1010011000001000000000000000", -- 336                                                       jump      _42
"1010101011000000000000001110", -- 337 alu-gc              free                              num?      _46
"0000000000000000000101001110", -- 338 _45                 free       mar                    
"0000000000000000000110100010", -- 339                     mem        free                   
"0000000001101000000000100100", -- 340                     buf1       bidir                  return    
"1010101111100000000000000000", -- 341 _46                                                   call      gc
"1010100100001000000000000000", -- 342                                                       jump      _45
"1011011111100100100111100111", -- 343 gc                  s          root       gc          call      mark-start
"1011011111100000000111101000", -- 344                     e          root                   call      mark-start
"1011011111100000000111101001", -- 345                     c          root                   call      mark-start
"1011011111100000000111101010", -- 346                     d          root                   call      mark-start
"1011011111100000000111101100", -- 347                     x1         root                   call      mark-start
"1011011111100000000111101101", -- 348                     x2         root                   call      mark-start
"1011011111100000000111110100", -- 349                     nilx       root                   call      mark-start
"1011011111100000000111110101", -- 350                     true       root                   call      mark-start
"1011011111100000000111110110", -- 351                     false      root                   call      mark-start
"0000000000000000000110110011", -- 352                     num        free                   
"0000000000000000000001010011", -- 353                     num        arg                    
"0000000000000000010010000000", -- 354                                buf2       dec         
"0000000000000000000101000101", -- 355                     buf2       mar                    
"1011011011010000000000000011", -- 356 _48                 arg                               nil?      _51
"1011010000011000000001000010", -- 357                     mem        arg                    mark?     _49
"0000000000000000000000101110", -- 358                     free       bidir                  
"1011010100001000000110101011", -- 359                     mar        free                   jump      _50
"0000000000000010010010000000", -- 360 _49                            buf2       clear-mark  
"0000000000000000000000100101", -- 361                     buf2       bidir                  
"0000000000000000000001001011", -- 362 _50                 mar        arg                    
"0000000000000000010010000000", -- 363                                buf2       dec         
"1011001000001000000101000101", -- 364                     buf2       mar                    jump      _48
"0000110011000000000000001110", -- 365 _51                 free                              num?      error
"0000000001101100000000000000", -- 366                                           running     return    
"0000000000000000000111010100", -- 367 mark-start          nilx       parent                 
"0000000000000000000101010000", -- 368 mark                root       mar                    
"1011110000011000000001000010", -- 369                     mem        arg                    mark?     backup
"0000000000000001110010000000", -- 370                                buf2       set-mark    
"1011110001001000000000100101", -- 371                     buf2       bidir                  atom?     backup
"0000000000000000001000001111", -- 372                     parent     y1                     
"0000000000000000001000110000", -- 373                     root       y2                     
"0000000000000011110000000000", -- 374                                           gcmark      
"1011100000001000000000100101", -- 375                     buf2       bidir                  jump      mark
"1100000011010000000101001111", -- 376 backup              parent     mar                    nil?      _56
"1011111100100000000001000010", -- 377                     mem        arg                    field?    _55
"0000000000000000001000010000", -- 378                     root       y1                     
"0000000000000000001000101111", -- 379                     parent     y2                     
"0000000000000011100000000000", -- 380                                           gcreset     
"1011110000001000000000100101", -- 381                     buf2       bidir                  jump      backup
"0000000000000000001000110000", -- 382 _55                 root       y2                     
"0000000000000011010000000000", -- 383                                           gcreverse   
"1011100000001000000000100101", -- 384                     buf2       bidir                  jump      mark
"0000000001101000000000000000", -- 385 _56                                                   return    
others => (others => '0'));

begin

  process (clk)
  begin
    if falling_edge(clk) then
      if en = '1' then
        data <= MICROCODE_ROM(conv_integer(addr));
      end if;
    end if;
  end process;


end;

