

-- Automatically generated SECD microcode

library ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity microcode_rom is
  port (clk  : in std_logic;
        en   : in std_logic;
        addr : in std_logic_vector(8 downto 0);
        data : out std_logic_vector(27 downto 0));
end microcode_rom;

architecture rtl of microcode_rom is

constant MICROCODE_ROM_SIZE : integer := 512;
type rom_type is array (0 to MICROCODE_ROM_SIZE - 1) of std_logic_vector (27 downto 0);
constant MICROCODE_ROM : rom_type := (
"0001001000001000000000000000", -- 0                                                         jump      boot
"0001111100001000000000000000", -- 1   ld-ins                                                jump      ld
"0011001010001000000000000000", -- 2   ldc-ins                                               jump      ldc
"0011100000001000000000000000", -- 3   ldf-ins                                               jump      ldf
"0011111010001000000000000000", -- 4   ap-ins                                                jump      ap
"0100110010001000000000000000", -- 5   rtn-ins                                               jump      rtn
"0101011000001000000000000000", -- 6   dum-ins                                               jump      dum
"0101100010001000000000000000", -- 7   rap-ins                                               jump      rap
"0110100000001000000000000000", -- 8   sel-ins                                               jump      sel
"0111011000001000000000000000", -- 9   join-ins                                              jump      join
"1000101100001000000000000000", -- 10  car-ins                                               jump      car
"1001000000001000000000000000", -- 11  cdr-ins                                               jump      cdr
"1001010010001000000000000000", -- 12  atom-ins                                              jump      atom
"1001101000001000000000000000", -- 13  cons-ins                                              jump      cons
"1010001000001000000000000000", -- 14  eq-ins                                                jump      eq
"1010010100001000000000000000", -- 15  add-ins                                               jump      add
"1010011100001000000000000000", -- 16  sub-ins                                               jump      sub
"1010100100001000000000000000", -- 17  mul-ins                                               jump      mul
"1010101100001000000000000000", -- 18  div-ins                                               jump      div
"1010110100001000000000000000", -- 19  rem-ins                                               jump      rem
"1010111100001000000000000000", -- 20  leq-ins                                               jump      leq
"1011001000001000000000000000", -- 21  stop-ins                                              jump      stop
"1011010010001000000000000000", -- 22  external-ins                                          jump      external
"1011001000001000000000000000", -- 23  cmd23-ins                                             jump      stop
"1011001000001000000000000000", -- 24  cmd24-ins                                             jump      stop
"1011001000001000000000000000", -- 25  cmd25-ins                                             jump      stop
"1011001000001000000000000000", -- 26  cmd26-ins                                             jump      stop
"1011001000001000000000000000", -- 27  cmd27-ins                                             jump      stop
"1011001000001000000000000000", -- 28  cmd28-ins                                             jump      stop
"1011001000001000000000000000", -- 29  cmd29-ins                                             jump      stop
"1011001000001000000000000000", -- 30  cmd30-ins                                             jump      stop
"0111100100001000000000000000", -- 31  fork-ins                                              jump      fork
"1000010010001000000000000000", -- 32  fail-ins                                              jump      fail
"1011001000001000000000000000", -- 33  delay-ins                                             jump      stop
"1011001000001000000000000000", -- 34  delay0-ins                                            jump      stop
"1011001000001000000000000000", -- 35  force-ins                                             jump      stop
"0001010101011100010000000000", -- 36  boot            1                         halted      button?   start-program
"0001001000001000000000000000", -- 37                                                        jump      boot
"0001010001011000000000000000", -- 38  error           2                                     button?   _3
"0001001100001000000000000000", -- 39                                                        jump      error
"0001010001011000000000000000", -- 40  _3                                                    button?   _3
"0001001000001000000000000000", -- 41                                                        jump      boot
"0000000000000100000101010011", -- 42  start-program       num        mar        running     
"0000000000000000000010100010", -- 43                      mem        car                    
"0000000000000000000101000110", -- 44                      car        mar                    
"0000000000000000000011000010", -- 45                      mem        s                      
"0000000000000000000011110100", -- 46                      nilx       e                      
"0000000000000000000101010011", -- 47                      num        mar                    
"0000000000000000000010100010", -- 48                      mem        car                    
"0000000000000000000101000110", -- 49                      car        mar                    
"0000000000000000000010100010", -- 50                      mem        car                    
"0000000000000000000100000110", -- 51                      car        c                      
"0000000000000000000100110100", -- 52                      nilx       d                      
"0000000000000000000101110100", -- 53                      nilx       x1                     
"0000000000000000000110010100", -- 54                      nilx       x2                     
"0000000000000000001001010100", -- 55                      nilx       r                      
"0000000000000000000101010011", -- 56                      num        mar                    
"0000000000000000000110100010", -- 57                      mem        free                   
"0000000000000000000101001001", -- 58  top-of-cycle        c          mar                    
"0000000000000000000010100010", -- 59                      mem        car                    
"0000000000000000000101000110", -- 60                      car        mar                    
"0000000000010000000001000010", -- 61                      mem        arg                    dispatch  
"0000000000000000000101101000", -- 62  ld                  e          x1                     
"0000000000000000000101001001", -- 63                      c          mar                    
"0000000000000000000110000010", -- 64                      mem        x2                     
"0000000000000000000101001101", -- 65                      x2         mar                    
"0000000000000000000010100010", -- 66                      mem        car                    
"0000000000000000000101000110", -- 67                      car        mar                    
"0000000000000000000010100010", -- 68                      mem        car                    
"0000000000000000000101000110", -- 69                      car        mar                    
"0000000000000000000001000010", -- 70                      mem        arg                    
"0010011001010000000000000011", -- 71  _7                  arg                               nil?      _8
"0000000000000000000101001100", -- 72                      x1         mar                    
"0000000000000000000101100010", -- 73                      mem        x1                     
"0000000000000000010001100000", -- 74                                 buf1       dec         
"0010001110001000000001000100", -- 75                      buf1       arg                    jump      _7
"0000000000000000000101001100", -- 76  _8                  x1         mar                    
"0000000000000000000010100010", -- 77                      mem        car                    
"0000000000000000000101100110", -- 78                      car        x1                     
"0000000000000000000101001001", -- 79                      c          mar                    
"0000000000000000000110000010", -- 80                      mem        x2                     
"0000000000000000000101001101", -- 81                      x2         mar                    
"0000000000000000000010100010", -- 82                      mem        car                    
"0000000000000000000101000110", -- 83                      car        mar                    
"0000000000000000000110000010", -- 84                      mem        x2                     
"0000000000000000000101001101", -- 85                      x2         mar                    
"0000000000000000000001000010", -- 86                      mem        arg                    
"0010111001010000000000000011", -- 87  _9                  arg                               nil?      _10
"0000000000000000000101001100", -- 88                      x1         mar                    
"0000000000000000000101100010", -- 89                      mem        x1                     
"0000000000000000010001100000", -- 90                                 buf1       dec         
"0010101110001000000001000100", -- 91                      buf1       arg                    jump      _9
"0000000000000000000101001100", -- 92  _10                 x1         mar                    
"0000000000000000000010100010", -- 93                      mem        car                    
"0000000000000000000101100110", -- 94                      car        x1                     
"1011111011100000000110000111", -- 95                      s          x2                     call      consx1x2
"0000000000000000000011001011", -- 96                      mar        s                      
"0000000000000000000101001001", -- 97                      c          mar                    
"0000000000000000000100000010", -- 98                      mem        c                      
"0000000000000000000101001001", -- 99                      c          mar                    
"0001110100001000000100000010", -- 100                     mem        c                      jump      top-of-cycle
"0000000000000000000110000111", -- 101 ldc                 s          x2                     
"0000000000000000000101001001", -- 102                     c          mar                    
"0000000000000000000101100010", -- 103                     mem        x1                     
"0000000000000000000101001100", -- 104                     x1         mar                    
"0000000000000000000010100010", -- 105                     mem        car                    
"1011111011100000000101100110", -- 106                     car        x1                     call      consx1x2
"0000000000000000000011001011", -- 107                     mar        s                      
"0000000000000000000101001001", -- 108                     c          mar                    
"0000000000000000000100000010", -- 109                     mem        c                      
"0000000000000000000101001001", -- 110                     c          mar                    
"0001110100001000000100000010", -- 111                     mem        c                      jump      top-of-cycle
"0000000000000000000110001000", -- 112 ldf                 e          x2                     
"0000000000000000000101001001", -- 113                     c          mar                    
"0000000000000000000101100010", -- 114                     mem        x1                     
"0000000000000000000101001100", -- 115                     x1         mar                    
"0000000000000000000010100010", -- 116                     mem        car                    
"1011111011100000000101100110", -- 117                     car        x1                     call      consx1x2
"0000000000000000000101101011", -- 118                     mar        x1                     
"1011111011100000000110000111", -- 119                     s          x2                     call      consx1x2
"0000000000000000000011001011", -- 120                     mar        s                      
"0000000000000000000101001001", -- 121                     c          mar                    
"0000000000000000000100000010", -- 122                     mem        c                      
"0000000000000000000101001001", -- 123                     c          mar                    
"0001110100001000000100000010", -- 124                     mem        c                      jump      top-of-cycle
"0000000000000000000110001010", -- 125 ap                  d          x2                     
"0000000000000000000101001001", -- 126                     c          mar                    
"1011111011100000000101100010", -- 127                     mem        x1                     call      consx1x2
"0000000000000000000110001011", -- 128                     mar        x2                     
"1011111011100000000101101000", -- 129                     e          x1                     call      consx1x2
"0000000000000000000110001011", -- 130                     mar        x2                     
"0000000000000000000101000111", -- 131                     s          mar                    
"0000000000000000000101100010", -- 132                     mem        x1                     
"0000000000000000000101001100", -- 133                     x1         mar                    
"1011111011100000000101100010", -- 134                     mem        x1                     call      consx1x2
"0000000000000000000100101011", -- 135                     mar        d                      
"0000000000000000000101000111", -- 136                     s          mar                    
"0000000000000000000010100010", -- 137                     mem        car                    
"0000000000000000000101000110", -- 138                     car        mar                    
"0000000000000000000110000010", -- 139                     mem        x2                     
"0000000000000000000101000111", -- 140                     s          mar                    
"0000000000000000000101100010", -- 141                     mem        x1                     
"0000000000000000000101001100", -- 142                     x1         mar                    
"0000000000000000000010100010", -- 143                     mem        car                    
"1011111011100000000101100110", -- 144                     car        x1                     call      consx1x2
"0000000000000000000011101011", -- 145                     mar        e                      
"0000000000000000000000000000", -- 146                                                       
"0000000000000000000101000111", -- 147                     s          mar                    
"0000000000000000000010100010", -- 148                     mem        car                    
"0000000000000000000101000110", -- 149                     car        mar                    
"0000000000000000000010100010", -- 150                     mem        car                    
"0000000000000000000100000110", -- 151                     car        c                      
"0001110100001000000011010100", -- 152                     nilx       s                      jump      top-of-cycle
"0000000000000000000101001010", -- 153 rtn                 d          mar                    
"0000000000000000000010100010", -- 154                     mem        car                    
"0000000000000000000110000110", -- 155                     car        x2                     
"0000000000000000000101000111", -- 156                     s          mar                    
"0000000000000000000010100010", -- 157                     mem        car                    
"1011111011100000000101100110", -- 158                     car        x1                     call      consx1x2
"0000000000000000000011001011", -- 159                     mar        s                      
"0000000000000000000101001010", -- 160                     d          mar                    
"0000000000000000000100100010", -- 161                     mem        d                      
"0000000000000000000101001010", -- 162                     d          mar                    
"0000000000000000000010100010", -- 163                     mem        car                    
"0000000000000000000011100110", -- 164                     car        e                      
"0000000000000000000101001010", -- 165                     d          mar                    
"0000000000000000000100100010", -- 166                     mem        d                      
"0000000000000000000101001010", -- 167                     d          mar                    
"0000000000000000000010100010", -- 168                     mem        car                    
"0000000000000000000100000110", -- 169                     car        c                      
"0000000000000000000101001010", -- 170                     d          mar                    
"0001110100001000000100100010", -- 171                     mem        d                      jump      top-of-cycle
"0000000000000000000110001000", -- 172 dum                 e          x2                     
"1011111011100000000101110100", -- 173                     nilx       x1                     call      consx1x2
"0000000000000000000011101011", -- 174                     mar        e                      
"0000000000000000000101001001", -- 175                     c          mar                    
"0001110100001000000100000010", -- 176                     mem        c                      jump      top-of-cycle
"0000000000000000000110001010", -- 177 rap                 d          x2                     
"0000000000000000000101001001", -- 178                     c          mar                    
"1011111011100000000101100010", -- 179                     mem        x1                     call      consx1x2
"0000000000000000000110001011", -- 180                     mar        x2                     
"0000000000000000000101001000", -- 181                     e          mar                    
"1011111011100000000101100010", -- 182                     mem        x1                     call      consx1x2
"0000000000000000000110001011", -- 183                     mar        x2                     
"0000000000000000000101000111", -- 184                     s          mar                    
"0000000000000000000101100010", -- 185                     mem        x1                     
"0000000000000000000101001100", -- 186                     x1         mar                    
"1011111011100000000101100010", -- 187                     mem        x1                     call      consx1x2
"0000000000000000000100101011", -- 188                     mar        d                      
"0000000000000000000101000111", -- 189                     s          mar                    
"0000000000000000000010100010", -- 190                     mem        car                    
"0000000000000000000101000110", -- 191                     car        mar                    
"0000000000000000000011100010", -- 192                     mem        e                      
"0000000000000000000101000111", -- 193                     s          mar                    
"0000000000000000001000100010", -- 194                     mem        y2                     
"0000000000000000000101010010", -- 195                     y2         mar                    
"0000000000000000000010100010", -- 196                     mem        car                    
"0000000000000000001000100110", -- 197                     car        y2                     
"0000000000000000000101001000", -- 198                     e          mar                    
"0000000000000000000001000010", -- 199                     mem        arg                    
"0000000000000010100001100000", -- 200                                buf1       replcar     
"0000000000000000000000100100", -- 201                     buf1       bidir                  
"0000000000000000000101000111", -- 202                     s          mar                    
"0000000000000000000010100010", -- 203                     mem        car                    
"0000000000000000000101000110", -- 204                     car        mar                    
"0000000000000000000010100010", -- 205                     mem        car                    
"0000000000000000000100000110", -- 206                     car        c                      
"0001110100001000000011010100", -- 207                     nilx       s                      jump      top-of-cycle
"0000000000000000000110001010", -- 208 sel                 d          x2                     
"0000000000000000000101001001", -- 209                     c          mar                    
"0000000000000000000101100010", -- 210                     mem        x1                     
"0000000000000000000101001100", -- 211                     x1         mar                    
"0000000000000000000101100010", -- 212                     mem        x1                     
"0000000000000000000101001100", -- 213                     x1         mar                    
"1011111011100000000101100010", -- 214                     mem        x1                     call      consx1x2
"0000000000000000000100101011", -- 215                     mar        d                      
"0000000000000000000101000111", -- 216                     s          mar                    
"0000000000000000000010100010", -- 217                     mem        car                    
"0000000000000000000101000110", -- 218                     car        mar                    
"0000000000000000000001000010", -- 219                     mem        arg                    
"0000000000000000000101010101", -- 220                     true       mar                    
"0111001010110000000000000010", -- 221                     mem                               eq?       _18
"0000000000000000000101001001", -- 222                     c          mar                    
"0000000000000000000100000010", -- 223                     mem        c                      
"0000000000000000000101001001", -- 224                     c          mar                    
"0000000000000000000100000010", -- 225                     mem        c                      
"0000000000000000000101001001", -- 226                     c          mar                    
"0000000000000000000010100010", -- 227                     mem        car                    
"0111010100001000000100000110", -- 228                     car        c                      jump      _19
"0000000000000000000101001001", -- 229 _18                 c          mar                    
"0000000000000000000100000010", -- 230                     mem        c                      
"0000000000000000000101001001", -- 231                     c          mar                    
"0000000000000000000010100010", -- 232                     mem        car                    
"0000000000000000000100000110", -- 233                     car        c                      
"0000000000000000000101000111", -- 234 _19                 s          mar                    
"0001110100001000000011000010", -- 235                     mem        s                      jump      top-of-cycle
"0000000000000000000100001010", -- 236 join                d          c                      
"0000000000000000000101001001", -- 237                     c          mar                    
"0000000000000000000010100010", -- 238                     mem        car                    
"0000000000000000000100000110", -- 239                     car        c                      
"0000000000000000000101001010", -- 240                     d          mar                    
"0001110100001000000100100010", -- 241                     mem        d                      jump      top-of-cycle
"0000000000000000000101001001", -- 242 fork                c          mar                    
"0000000000000000000101000010", -- 243                     mem        mar                    
"0000000000000000000101000010", -- 244                     mem        mar                    
"0000000000000000000101100010", -- 245                     mem        x1                     
"1011111011100000000110001010", -- 246                     d          x2                     call      consx1x2
"0000000000000000000100101011", -- 247                     mar        d                      
"0000000000000000000101101011", -- 248                     mar        x1                     
"1011111011100000000110011000", -- 249                     r          x2                     call      consx1x2
"0000000000000000000110001011", -- 250                     mar        x2                     
"0000000000000000000101001001", -- 251                     c          mar                    
"0000000000000000000101000010", -- 252                     mem        mar                    
"0000000000000000000101000010", -- 253                     mem        mar                    
"0000000000000000000010100010", -- 254                     mem        car                    
"1011111011100000000101100110", -- 255                     car        x1                     call      consx1x2
"0000000000000000000110001011", -- 256                     mar        x2                     
"1011111011100000000101101000", -- 257                     e          x1                     call      consx1x2
"0000000000000000000110001011", -- 258                     mar        x2                     
"1011111011100000000101100111", -- 259                     s          x1                     call      consx1x2
"0000000000000000001001001011", -- 260                     mar        r                      
"0000000000000000000101001001", -- 261                     c          mar                    
"0000000000000000000101000010", -- 262                     mem        mar                    
"0000000000000000000010100010", -- 263                     mem        car                    
"0001110100001000000100000110", -- 264                     car        c                      jump      top-of-cycle
"0000000000000000000101011000", -- 265 fail                r          mar                    
"0000000000000000000010100010", -- 266                     mem        car                    
"0000000000000000000011000110", -- 267                     car        s                      
"0000000000000000000101000010", -- 268                     mem        mar                    
"0000000000000000000010100010", -- 269                     mem        car                    
"0000000000000000000011100110", -- 270                     car        e                      
"0000000000000000000101000010", -- 271                     mem        mar                    
"0000000000000000000010100010", -- 272                     mem        car                    
"0000000000000000000100000110", -- 273                     car        c                      
"0000000000000000000101000010", -- 274                     mem        mar                    
"0000000000000000000010100010", -- 275                     mem        car                    
"0000000000000000000100100110", -- 276                     car        d                      
"0001110100001000001001000010", -- 277                     mem        r                      jump      top-of-cycle
"0000000000000000000101000111", -- 278 car                 s          mar                    
"0000000000000000000110000010", -- 279                     mem        x2                     
"0000000000000000000101000111", -- 280                     s          mar                    
"0000000000000000000010100010", -- 281                     mem        car                    
"0000000000000000000101000110", -- 282                     car        mar                    
"0000000000000000000010100010", -- 283                     mem        car                    
"1011111011100000000101100110", -- 284                     car        x1                     call      consx1x2
"0000000000000000000011001011", -- 285                     mar        s                      
"0000000000000000000101001001", -- 286                     c          mar                    
"0001110100001000000100000010", -- 287                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 288 cdr                 s          mar                    
"0000000000000000000110000010", -- 289                     mem        x2                     
"0000000000000000000101000111", -- 290                     s          mar                    
"0000000000000000000010100010", -- 291                     mem        car                    
"0000000000000000000101000110", -- 292                     car        mar                    
"1011111011100000000101100010", -- 293                     mem        x1                     call      consx1x2
"0000000000000000000011001011", -- 294                     mar        s                      
"0000000000000000000101001001", -- 295                     c          mar                    
"0001110100001000000100000010", -- 296                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 297 atom                s          mar                    
"0000000000000000000010100010", -- 298                     mem        car                    
"0000000000000000000101000110", -- 299                     car        mar                    
"1001011101001000000000000010", -- 300                     mem                               atom?     _24
"1001011110001000000101110110", -- 301                     false      x1                     jump      _25
"0000000000000000000101110101", -- 302 _24                 true       x1                     
"0000000000000000000101000111", -- 303 _25                 s          mar                    
"1011111011100000000110000010", -- 304                     mem        x2                     call      consx1x2
"0000000000000000000011001011", -- 305                     mar        s                      
"0000000000000000000101001001", -- 306                     c          mar                    
"0001110100001000000100000010", -- 307                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 308 cons                s          mar                    
"0000000000000000000110000010", -- 309                     mem        x2                     
"0000000000000000000101001101", -- 310                     x2         mar                    
"0000000000000000000010100010", -- 311                     mem        car                    
"0000000000000000000110000110", -- 312                     car        x2                     
"0000000000000000000101000111", -- 313                     s          mar                    
"0000000000000000000010100010", -- 314                     mem        car                    
"1011111011100000000101100110", -- 315                     car        x1                     call      consx1x2
"0000000000000000000101101011", -- 316                     mar        x1                     
"0000000000000000000101000111", -- 317                     s          mar                    
"0000000000000000000110000010", -- 318                     mem        x2                     
"0000000000000000000101001101", -- 319                     x2         mar                    
"1011111011100000000110000010", -- 320                     mem        x2                     call      consx1x2
"0000000000000000000011001011", -- 321                     mar        s                      
"0000000000000000000101001001", -- 322                     c          mar                    
"0001110100001000000100000010", -- 323                     mem        c                      jump      top-of-cycle
"1011011011100000000000000000", -- 324 eq                                                    call      setup-alu-args
"1010001110110000000000000010", -- 325                     mem                               eq?       _28
"1010010000001000000101110110", -- 326                     false      x1                     jump      _29
"0000000000000000000101110101", -- 327 _28                 true       x1                     
"1011101101100000000000000000", -- 328 _29                                                   call      push-alu-result
"0001110100001000000000000000", -- 329                                                       jump      top-of-cycle
"1011011011100000000000000000", -- 330 add                                                   call      setup-alu-args
"1100000111100000100001100010", -- 331                     mem        buf1       add         call      alu-gc
"1011101101100000000101101011", -- 332                     mar        x1                     call      push-alu-result
"0001110100001000000000000000", -- 333                                                       jump      top-of-cycle
"1011011011100000000000000000", -- 334 sub                                                   call      setup-alu-args
"1100000111100000110001100010", -- 335                     mem        buf1       sub         call      alu-gc
"1011101101100000000101101011", -- 336                     mar        x1                     call      push-alu-result
"0001110100001000000000000000", -- 337                                                       jump      top-of-cycle
"1011011011100000000000000000", -- 338 mul                                                   call      setup-alu-args
"1100000111100001000001100010", -- 339                     mem        buf1       mul         call      alu-gc
"1011101101100000000101101011", -- 340                     mar        x1                     call      push-alu-result
"0001110100001000000000000000", -- 341                                                       jump      top-of-cycle
"1011011011100000000000000000", -- 342 div                                                   call      setup-alu-args
"1100000111100001010001100010", -- 343                     mem        buf1       div         call      alu-gc
"1011101101100000000101101011", -- 344                     mar        x1                     call      push-alu-result
"0001110100001000000000000000", -- 345                                                       jump      top-of-cycle
"1011011011100000000000000000", -- 346 rem                                                   call      setup-alu-args
"1100000111100001100001100010", -- 347                     mem        buf1       rem         call      alu-gc
"1011101101100000000101101011", -- 348                     mar        x1                     call      push-alu-result
"0001110100001000000000000000", -- 349                                                       jump      top-of-cycle
"1011011011100000000000000000", -- 350 leq                                                   call      setup-alu-args
"1011000010111000000000000010", -- 351                     mem                               leq?      _36
"1011000100001000000101110110", -- 352                     false      x1                     jump      _37
"0000000000000000000101110101", -- 353 _36                 true       x1                     
"1011101101100000000000000000", -- 354 _37                                                   call      push-alu-result
"0001110100001000000000000000", -- 355                                                       jump      top-of-cycle
"0000000000000000000101000111", -- 356 stop                s          mar                    
"0000000000000000000010100010", -- 357                     mem        car                    
"0000000000000000000011000110", -- 358                     car        s                      
"0000000000000000000101010011", -- 359                     num        mar                    
"0000000001110000000000100111", -- 360                     s          bidir                  stop      
"1011010111011100110000000000", -- 361 external                                  external    button?   external-finish
"1011010010001000000000000000", -- 362                                                       jump      external
"0000000000000100000101001001", -- 363 external-finish     c          mar        running     
"0001110100001000000100000010", -- 364                     mem        c                      jump      top-of-cycle
"0000000000000000000101000111", -- 365 setup-alu-args      s          mar                    
"0000000000000000000101100010", -- 366                     mem        x1                     
"0000000000000000000101001100", -- 367                     x1         mar                    
"0000000000000000000010100010", -- 368                     mem        car                    
"0000000000000000000101000110", -- 369                     car        mar                    
"0000000000000000000001000010", -- 370                     mem        arg                    
"0000000000000000000101000111", -- 371                     s          mar                    
"0000000000000000000010100010", -- 372                     mem        car                    
"0000000001101000000101000110", -- 373                     car        mar                    return    
"0000000000000000000101000111", -- 374 push-alu-result     s          mar                    
"0000000000000000000110000010", -- 375                     mem        x2                     
"0000000000000000000101001101", -- 376                     x2         mar                    
"1011111011100000000110000010", -- 377                     mem        x2                     call      consx1x2
"0000000000000000000011001011", -- 378                     mar        s                      
"0000000000000000000101001001", -- 379                     c          mar                    
"0000000001101000000100000010", -- 380                     mem        c                      return    
"1100000011000000000000001110", -- 381 consx1x2            free                              num?      cons-gc
"0000000000000000000101001110", -- 382 _42                 free       mar                    
"0000000000000000000110100010", -- 383                     mem        free                   
"0000000001101000000000110111", -- 384                     cons       bidir                  return    
"1100010011100000000000000000", -- 385 cons-gc                                               call      gc
"1011111100001000000000000000", -- 386                                                       jump      _42
"1100001111000000000000001110", -- 387 alu-gc              free                              num?      _46
"0000000000000000000101001110", -- 388 _45                 free       mar                    
"0000000000000000000110100010", -- 389                     mem        free                   
"0000000001101000000000100100", -- 390                     buf1       bidir                  return    
"1100010011100000000000000000", -- 391 _46                                                   call      gc
"1100001000001000000000000000", -- 392                                                       jump      _45
"1101000101100100100111100111", -- 393 gc                  s          root       gc          call      mark-start
"1101000101100000000111101000", -- 394                     e          root                   call      mark-start
"1101000101100000000111101001", -- 395                     c          root                   call      mark-start
"1101000101100000000111101010", -- 396                     d          root                   call      mark-start
"1101000101100000000111111000", -- 397                     r          root                   call      mark-start
"1101000101100000000111101100", -- 398                     x1         root                   call      mark-start
"1101000101100000000111101101", -- 399                     x2         root                   call      mark-start
"1101000101100000000111110100", -- 400                     nilx       root                   call      mark-start
"1101000101100000000111110101", -- 401                     true       root                   call      mark-start
"1101000101100000000111110110", -- 402                     false      root                   call      mark-start
"0000000000000000000110110011", -- 403                     num        free                   
"0000000000000000000001010011", -- 404                     num        arg                    
"0000000000000000010010000000", -- 405                                buf2       dec         
"0000000000000000000101000101", -- 406                     buf2       mar                    
"1101000001010000000000000011", -- 407 _48                 arg                               nil?      _51
"1100110110011000000001000010", -- 408                     mem        arg                    mark?     _49
"0000000000000000000000101110", -- 409                     free       bidir                  
"1100111010001000000110101011", -- 410                     mar        free                   jump      _50
"0000000000000010010010000000", -- 411 _49                            buf2       clear-mark  
"0000000000000000000000100101", -- 412                     buf2       bidir                  
"0000000000000000000001001011", -- 413 _50                 mar        arg                    
"0000000000000000010010000000", -- 414                                buf2       dec         
"1100101110001000000101000101", -- 415                     buf2       mar                    jump      _48
"0001001101000000000000001110", -- 416 _51                 free                              num?      error
"0000000001101100000000000000", -- 417                                           running     return    
"0000000000000000000111010100", -- 418 mark-start          nilx       parent                 
"0000000000000000000101010000", -- 419 mark                root       mar                    
"1101010110011000000001000010", -- 420                     mem        arg                    mark?     backup
"0000000000000001110010000000", -- 421                                buf2       set-mark    
"1101010111001000000000100101", -- 422                     buf2       bidir                  atom?     backup
"0000000000000000001000001111", -- 423                     parent     y1                     
"0000000000000000001000110000", -- 424                     root       y2                     
"0000000000000011110000000000", -- 425                                           gcmark      
"1101000110001000000000100101", -- 426                     buf2       bidir                  jump      mark
"1101101001010000000101001111", -- 427 backup              parent     mar                    nil?      _56
"1101100010100000000001000010", -- 428                     mem        arg                    field?    _55
"0000000000000000001000010000", -- 429                     root       y1                     
"0000000000000000001000101111", -- 430                     parent     y2                     
"0000000000000011100000000000", -- 431                                           gcreset     
"1101010110001000000000100101", -- 432                     buf2       bidir                  jump      backup
"0000000000000000001000110000", -- 433 _55                 root       y2                     
"0000000000000011010000000000", -- 434                                           gcreverse   
"1101000110001000000000100101", -- 435                     buf2       bidir                  jump      mark
"0000000001101000000000000000", -- 436 _56                                                   return    
others => (others => '0'));

begin

  process (clk)
  begin
    if falling_edge(clk) then
      if en = '1' then
        data <= MICROCODE_ROM(conv_integer(addr));
      end if;
    end if;
  end process;


end;

